library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Noisy_Signal_Generation is
     Port (
         clk                  : in  std_logic := '0';           -- Clock signal
         reset                : in  std_logic := '0';           -- Reset signal
         x_out                : Out signed(15 downto 0):= (others=>'0');   
         sample_valid_Out     : out std_logic := '0'      -- Sample valid input signal
     );
end Noisy_Signal_Generation;

architecture Behavioral of Noisy_Signal_Generation is
 
signal clockcounter : integer range 0 to 64; 

type InputData_Array is array(0 to 1559) of signed(15 downto 0);  -- need 27 bits
    signal InputData : InputData_Array := (  
    
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16)
); 

begin

process(clk,reset)
variable index: integer:= 0; 
begin
     if(reset='1') then
         clockcounter<=0;
         sample_valid_Out<='0';
     elsif(rising_edge(clk)) then
         clockcounter <=clockcounter+1;
             if (clockcounter=64) then
                 sample_valid_Out <='1'; 
                 clockcounter<=0; 
                 x_out <= InputData(index);
                 index:= index+1; 
                       if(index = 1560) then 
                         index :=0; 
                       end if;
             else
                 sample_valid_Out <='0'; 
             end if;
     end if; 
end process;


end behavioral; 